module EA (
input [9:0] hsync,
input [9:0] vsync,
output reg [23:0] rgb );


reg [0:159] sprite [0:47];


always @(*) begin 

sprite[0] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[1] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[2] =  160'b0000000000000000000000000000000000000000000000000000000000000000000001111111100000111000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[3] =  160'b0000000000000000000000000000000000000000000000000000000000000000000001100000000000111000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[4] =  160'b0000000000000000000000000000000000000000000000000000000000000000000001100000000001111100000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[5] =  160'b0000000000000000000000000000000000000000000000000000000000000000000001100000000001101100000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[6] =  160'b0000000000000000000000000000000000000000000000000000000000000000000001100000000001101110000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[7] =  160'b0000000000000000000000000000000000000000000000000000000000000000000001111111000011000110000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[8] =  160'b0000000000000000000000000000000000000000000000000000000000000000000001111111000011000110000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[9] =  160'b0000000000000000000000000000000000000000000000000000000000000000000001100000000011000111000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[10] =  160'b0000000000000000000000000000000000000000000000000000000000000000000001100000000111111111000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[11] =  160'b0000000000000000000000000000000000000000000000000000000000000000000001100000000111111111000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[12] =  160'b0000000000000000000000000000000000000000000000000000000000000000000001100000000100000001100000000000000000000000000000000000000000000000000000000000000000000000;
sprite[13] =  160'b0000000000000000000000000000000000000000000000000000000000000000000001100000001100000001100000000000000000000000000000000000000000000000000000000000000000000000;
sprite[14] =  160'b0000000000000000000000000000000000000000000000000000000000000000000001111111101100000001100000000000000000000000000000000000000000000000000000000000000000000000;
sprite[15] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[16] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[17] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[18] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[19] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[20] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[21] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[22] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[23] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[24] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[25] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[26] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[27] =  160'b0000000000001100000000000000110000000000000000000000110001100000000000000001100000000000000000000000000110000000000000000000000000000001100000000000000000000000;
sprite[28] =  160'b0011111111001100000000000000110000000000000000000000110001100000000000000001100000000000111000000000000110000000000000000000000000000001100000000000000000000000;
sprite[29] =  160'b0011000000001100000000000000110000000011000000000000000001100000000000000000000000000000111000000000000110000000000000000000000000000001100000000000000000000000;
sprite[30] =  160'b0011000000001100000000000000110000000011000000000000000001100000000000000000000000000001111000000000000110000000000000000000000000000001100000000000000000000000;
sprite[31] =  160'b0011000000001100000011100000110001101111110001001100110001100011000011110001100000000001101100000001110110000011110000110011000011000001100000111100001100110000;
sprite[32] =  160'b0011000000001100001111111000110011101111110001111100110001100111000111111001100000000011001100000111111110001111111000111111111111110001100011111110001111110000;
sprite[33] =  160'b0011111110001100011000011000110111000011000001100000110001101110001100001001100000000011000100000110001110001000011000111000111000110001100010000110001110000000;
sprite[34] =  160'b0011111110001100011000001100111110000011000001100000110001111100001100000001100000000011000110000100000110000000001000110000110000110001100000000011001100000000;
sprite[35] =  160'b0011000000001100011111111100111100000011000001000000110001111000001000000001100000000110000110001100000110000011111000110000110000110001100000111111001100000000;
sprite[36] =  160'b0011000000001100011111111000111100000011000001000000110001111000001000000001100000000111111110001100000110001111111000110000110000110001100001111111001100000000;
sprite[37] =  160'b0011000000001100011000000000110110000011000001000000110001101100001000000001100000000111111111001100000110001100001000110000110000110001100011000011001100000000;
sprite[38] =  160'b0011000000001100011000000000110011000011000001000000110001100110001100000001100000001100000011000110000110001000001000110000110000110001100011000011001100000000;
sprite[39] =  160'b0011000000001100001100001000110011100011000001000000110001100111001110011001100000001100000001100111001110001100111000110000110000110001100011001111001100000000;
sprite[40] =  160'b0011111111001100000111111000110001110011110001000000110001100011100111110001100000011100000001100011111110001111101000110000110000110001100001111011001100000000;
sprite[41] =  160'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[42] =  160'b0000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[43] =  160'b0000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[44] =  160'b0000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[45] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[46] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[47] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
end

wire signed [9:0] x_rel, y_rel;
assign x_rel = hsync - 560;
assign y_rel = vsync - 44;

    always @(*) begin
        if (x_rel >= -80 && x_rel < 80 && y_rel >= -24 && y_rel < 24) begin
            if (sprite[y_rel + 24][x_rel + 80]) begin
                rgb = 24'hFFFF00;
				end
				else begin 
				rgb = 24'h000000;
				end
			end
			else begin
			rgb =24'h000000;
		end
    end
endmodule
