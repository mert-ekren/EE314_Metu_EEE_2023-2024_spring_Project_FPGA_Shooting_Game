module score_name(
input [9:0] hsync,
input [9:0] vsync,
output reg [23:0] rgb );

reg [0:159] sprite [0:39];

always @(*) begin

sprite[0] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[1] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[2] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[3] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[4] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[5] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[6] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[7] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[8] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[9] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[10] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[11] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[12] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[13] =  160'b0000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[14] =  160'b0000000000000000000000000000000000000000000000000000001100011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[15] =  160'b0000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[16] =  160'b0000000000000000000000000000000000000000000000000000011000000000011110000011110000011011100001110000000000110000000000000000000000000000000000000000000000000000;
sprite[17] =  160'b0000000000000000000000000000000000000000000000000000011100000000111111000111111100011111100111111100000000110000000000000000000000000000000000000000000000000000;
sprite[18] =  160'b0000000000000000000000000000000000000000000000000000001111000001110001001100001100011100000100001100000000110000000000000000000000000000000000000000000000000000;
sprite[19] =  160'b0000000000000000000000000000000000000000000000000000000111110001100000001100000110011000001100000110000000000000000000000000000000000000000000000000000000000000;
sprite[20] =  160'b0000000000000000000000000000000000000000000000000000000001111001100000001000000110011000001111111110000000000000000000000000000000000000000000000000000000000000;
sprite[21] =  160'b0000000000000000000000000000000000000000000000000000000000011001100000001000000110011000001111111100000000000000000000000000000000000000000000000000000000000000;
sprite[22] =  160'b0000000000000000000000000000000000000000000000000000000000011001100000001000000110011000001100000000000000000000000000000000000000000000000000000000000000000000;
sprite[23] =  160'b0000000000000000000000000000000000000000000000000000000000011001100000001100000110011000001100000000000000000000000000000000000000000000000000000000000000000000;
sprite[24] =  160'b0000000000000000000000000000000000000000000000000000011000111000110011001110011100011000000110000100000000110000000000000000000000000000000000000000000000000000;
sprite[25] =  160'b0000000000000000000000000000000000000000000000000000011111110000111111000111111000011000000011111100000000110000000000000000000000000000000000000000000000000000;
sprite[26] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[27] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[28] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[29] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[30] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[31] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[32] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[33] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[34] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[35] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[36] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[37] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[38] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[39] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;



end







wire signed [9:0] x_rel, y_rel;
assign x_rel = hsync - 560;
assign y_rel = vsync - 130;

    always @(*) begin
        if (x_rel >= -80 && x_rel < 80 && y_rel >= -20 && y_rel < 20) begin
            if (sprite[y_rel + 20][x_rel + 80]) begin
                rgb = 24'hFFFF00;
				end
				else begin 
				rgb = 24'h000000;
				end
			end
			else begin
			rgb =24'h000000;
		end
    end
endmodule

