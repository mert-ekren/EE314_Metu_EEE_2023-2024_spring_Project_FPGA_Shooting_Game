module over_drawing(
input[9:0]hcount,
input[9:0]vcount,
input reset,
input over,
output reg [23:0] rgb);

reg [0:127] sprite [0:31];
always @(*) begin

sprite[0] =  128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[1] =  128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[2] =  128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[3] =  128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[4] =  128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[5] =  128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[6] =  128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[7] =  128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[8] =  128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[9] =  128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[10] =  128'b00000000000000000000000000000000000001000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000;
sprite[11] =  128'b00000000001111100000000000000000000001000000000000001111111001000000000000000000000000000000000000000000000000000000000000000000;
sprite[12] =  128'b00000000001100110000000001100000000001000000000000000001100001000000000000000000000000000000000000000000000000000000000000000000;
sprite[13] =  128'b00000000001100110000000001100000000001000000000000000001100001000000000000000000000000000000000000000000000000000000000000000000;
sprite[14] =  128'b00000000001100110011110011110011110001001001111100000001100001111100011110000001111001111100010001001111011110011111000000000000;
sprite[15] =  128'b00000000001111100110001001100000011001010001000100000001100001000100110011000001000101000110010001001100010000010001000000000000;
sprite[16] =  128'b00000000001101100111111001100001111001100001111100000001100001000100111111000011000011000010010001001100011100011111000000000000;
sprite[17] =  128'b00000000001100100110000001100110011001010011000000000001100001000100100000000011000011000010010001001100000110110000000000000000;
sprite[18] =  128'b00000000001100110110000001100110011001011001000000000001100001000100110000000001000101000110010001001100000011010000000000000000;
sprite[19] =  128'b00000000001100010011111000110011111001001101111100000001100001000100011111000001111001111100011111001100011110011111000000000000;
sprite[20] =  128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[21] =  128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[22] =  128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[23] =  128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[24] =  128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[25] =  128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[26] =  128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[27] =  128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[28] =  128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[29] =  128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[30] =  128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[31] =  128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
end

wire signed [9:0] x_rel, y_rel;
assign x_rel = hcount - 240;
assign y_rel = vcount - 240;

    always @(*) begin
		if (reset) begin
		rgb =24'h000000;
		end
		else if (over) begin
        if (x_rel >= -64 && x_rel < 64 && y_rel >= -16 && y_rel < 16) begin
            if (sprite[y_rel + 16][x_rel + 64]) begin
                rgb = 24'hCC0066;
            end
				else begin 
				rgb =24'h202020;
				end
			end
			else begin
				rgb =24'h000000;
			end
		 end
		else begin
		rgb =24'h000000;
		end
    end
endmodule
