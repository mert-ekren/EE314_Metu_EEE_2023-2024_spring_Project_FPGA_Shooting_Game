module PlayerDrawing(
    input [3:0] angle_idx, // Angle index (0-15 for 0, 22.5, ..., 337.5 degrees)
    input [9:0] hcount, // Current horizontal pixel coordinate
    input [9:0] vcount, // Current vertical pixel coordinate
    input [9:0] x_center, // X coordinate of the player's center
    input [9:0] y_center, // Y coordinate of the player's center
    output reg [23:0] rgb // Output RGB value for the player pixel
);    
    // Define a 32x32 sprite
    reg [31:0] sprite [0:31];
    
    always @(*) begin
        case (angle_idx)
            4'd0: begin
                sprite[0] =  32'b00000000000000000000000000000000;
                sprite[1] =  32'b00000000000000000000000000000000;
                sprite[2] =  32'b00000000000000000000000000000000;
                sprite[3] =  32'b00000000000000000000000000000000;
                sprite[4] =  32'b00000000000000000000000000000000;
                sprite[5] =  32'b00000000000000001000000000000000;
                sprite[6] =  32'b00000000000000011100000000000000;
                sprite[7] =  32'b00000000000000111110000000000000;
                sprite[8] =  32'b00000000000000111110000000000000;
                sprite[9] =  32'b00000000000000111110000000000000;
                sprite[10] = 32'b00000000000001111111000000000000;
                sprite[11] = 32'b00000000000001111111000000000000;
                sprite[12] = 32'b00000000000001111111000000000000;
                sprite[13] = 32'b00000000000001111111000000000000;
                sprite[14] = 32'b00000000000011111111100000000000;
                sprite[15] = 32'b00000000000011111111100000000000;
                sprite[16] = 32'b00000000000011111111100000000000;
                sprite[17] = 32'b00000000000111111111110000000000;
                sprite[18] = 32'b00000000000111111111110000000000;
                sprite[19] = 32'b00000000000111111111110000000000;
                sprite[20] = 32'b00000000000111111111110000000000;
                sprite[21] = 32'b00000000000111111111110000000000;
                sprite[22] = 32'b00000000000111111111110000000000;
                sprite[23] = 32'b00000000000111111111110000000000;
                sprite[24] = 32'b00000000000000000000000000000000;
                sprite[25] = 32'b00000000000000000000000000000000;
                sprite[26] = 32'b00000000000000000000000000000000;
                sprite[27] = 32'b00000000000000000000000000000000;
                sprite[28] = 32'b00000000000000000000000000000000;
                sprite[29] = 32'b00000000000000000000000000000000;
                sprite[30] = 32'b00000000000000000000000000000000;
                sprite[31] = 32'b00000000000000000000000000000000;
            end 

				4'd1: begin
                sprite[0]  = 32'b00000000000000000000000000000000;
                sprite[1]  = 32'b00000000000000000000000000000000;
                sprite[2]  = 32'b00000000000000000000000000000000;
                sprite[3]  = 32'b00000000000000000000000000000000;
                sprite[4]  = 32'b00000000000000000000000000000000;
                sprite[5]  = 32'b00000000000000000000000000000000;
                sprite[6]  = 32'b00000000000000000000000000000000;
                sprite[7]  = 32'b00000000000000000000000000000000;
                sprite[8]  = 32'b00000000000000100000000000000000;
                sprite[9]  = 32'b00000000000011111000000000000000;
                sprite[10] = 32'b00000000000011111000000000000000;
                sprite[11] = 32'b00000000000011111110000000000000;
                sprite[12] = 32'b00000000000011111110000000000000;
                sprite[13] = 32'b00000000000001111110000000000000;
                sprite[14] = 32'b00000000000001111111110000000000;
                sprite[15] = 32'b00000000000000111111111000000000;
                sprite[16] = 32'b00000000000000111111111000000000;
                sprite[17] = 32'b00000000000000111111111110000000;
                sprite[18] = 32'b00000000000000111111111110000000;
                sprite[19] = 32'b00000000000000111111111110000000;
                sprite[20] = 32'b00000000000000011111111111000000;
                sprite[21] = 32'b00000000000000111111111100000000;
                sprite[22] = 32'b00000000000000111110000000000000;
                sprite[23] = 32'b00000000000000000000000000000000;
                sprite[24] = 32'b00000000000000000000000000000000;
                sprite[25] = 32'b00000000000000000000000000000000;
                sprite[26] = 32'b00000000000000000000000000000000;
                sprite[27] = 32'b00000000000000000000000000000000;
                sprite[28] = 32'b00000000000000000000000000000000;
                sprite[29] = 32'b00000000000000000000000000000000;
                sprite[30] = 32'b00000000000000000000000000000000;
                sprite[31] = 32'b00000000000000000000000000000000;
				end
				4'd2: begin
                sprite[0]  = 32'b00000000000000000000000000000000;
                sprite[1]  = 32'b00000000000000000000000000000000;
                sprite[2]  = 32'b00000000000000000000000000000000;
                sprite[3]  = 32'b00000000000000000000000000000000;
                sprite[4]  = 32'b00000000000000000000000000000000;
                sprite[5]  = 32'b00000000000000000000000000000000;
                sprite[6]  = 32'b00000000000000000000000000000000;
                sprite[7]  = 32'b00000000000000000000000000000000;
                sprite[8]  = 32'b00000000000000000000000000000000;
                sprite[9]  = 32'b00000000000000000000000000000000;
                sprite[10] = 32'b00000000000111000000000000000000;
                sprite[11] = 32'b00000000000111111100000000000000;
                sprite[12] = 32'b00000000000011111110000000000000;
                sprite[13] = 32'b00000000000001111111010000000000;
                sprite[14] = 32'b00000000000001111111111000000000;
                sprite[15] = 32'b00000000000001111111111110000000;
                sprite[16] = 32'b00000000000001111111111111000000;
                sprite[17] = 32'b00000000000000111111111111100000;
                sprite[18] = 32'b00000000000000011111111111100000;
                sprite[19] = 32'b00000000000000011111111111000000;
                sprite[20] = 32'b00000000000000001111111110000000;
                sprite[21] = 32'b00000000000000000111111100000000;
                sprite[22] = 32'b00000000000000001111111000000000;
                sprite[23] = 32'b00000000000000000111110000000000;
                sprite[24] = 32'b00000000000000000011100000000000;
                sprite[25] = 32'b00000000000000000000000000000000;
                sprite[26] = 32'b00000000000000000000000000000000;
                sprite[27] = 32'b00000000000000000000000000000000;
                sprite[28] = 32'b00000000000000000000000000000000;
                sprite[29] = 32'b00000000000000000000000000000000;
                sprite[30] = 32'b00000000000000000000000000000000;
                sprite[31] = 32'b00000000000000000000000000000000;
				end
				4'd3: begin
                sprite[0]  = 32'b00000000000000000000000000000000;
                sprite[1]  = 32'b00000000000000000000000000000000;
                sprite[2]  = 32'b00000000000000000000000000000000;
                sprite[3]  = 32'b00000000000000000000000000000000;
                sprite[4]  = 32'b00000000000000000000000000000000;
                sprite[5]  = 32'b00000000000000000000000000000000;
                sprite[6]  = 32'b00000000000000000000000000000000;
                sprite[7]  = 32'b00000000000000000000000000000000;
                sprite[8]  = 32'b00000000000000000000000000000000;
                sprite[9]  = 32'b00000000000000000000000000000000;
                sprite[10] = 32'b00000000000000000000000000000000;
                sprite[11] = 32'b00000000111111000000000000000000;
                sprite[12] = 32'b00000000111111111110000011100000;
                sprite[13] = 32'b00000000111111111111111110000000;
                sprite[14] = 32'b00000000111111111111111110000000;
                sprite[15] = 32'b00000000111111111111111100000000;
                sprite[16] = 32'b00000000000111111111111100000000;
                sprite[17] = 32'b00000000000111111111111000000000;
                sprite[18] = 32'b00000000000001111111111000000000;
                sprite[19] = 32'b00000000000000011111111110000000;
                sprite[20] = 32'b00000000000000001111111110000000;
                sprite[21] = 32'b00000000000000000011110000000000;
                sprite[22] = 32'b00000000000000000011100000000000;
                sprite[23] = 32'b00000000000000000001111000000000;
                sprite[24] = 32'b00000000000000000000000000000000;
                sprite[25] = 32'b00000000000000000000000000000000;
                sprite[26] = 32'b00000000000000000000000000000000;
                sprite[27] = 32'b00000000000000000000000000000000;
                sprite[28] = 32'b00000000000000000000000000000000;
                sprite[29] = 32'b00000000000000000000000000000000;
                sprite[30] = 32'b00000000000000000000000000000000;
                sprite[31] = 32'b00000000000000000000000000000000;
				end
					 4'd4: begin
                sprite[0]  = 32'b00000000000000000000000000000000;
                sprite[1]  = 32'b00000000000000000000000000000000;
                sprite[2]  = 32'b00000000000000000000000000000000;
                sprite[3]  = 32'b00000000000000000000000000000000;
                sprite[4]  = 32'b00000000000000000000000000000000;
                sprite[5]  = 32'b00000000000000000000000000000000;
                sprite[6]  = 32'b00000000000000000000000000000000;
                sprite[7]  = 32'b00000000000000000000000000000000;
                sprite[8]  = 32'b00000000000000000000000000000000;
                sprite[9]  = 32'b00000000000000000000000000000000;
                sprite[10] = 32'b00000000000000000000000000000000;
                sprite[11] = 32'b00000000000000111111110000000000;
                sprite[12] = 32'b00000000001111111111110000000000;
                sprite[13] = 32'b00000000111111111111110000000000;
                sprite[14] = 32'b00000011111111111111110000000000;
                sprite[15] = 32'b00000111111111111111110000000000;
                sprite[16] = 32'b00000011111111111111110000000000;
                sprite[17] = 32'b00000000111111111111110000000000;
                sprite[18] = 32'b00000000001111111111110000000000;
                sprite[19] = 32'b00000000000000111111110000000000;
                sprite[20] = 32'b00000000000000000000000000000000;
                sprite[21] = 32'b00000000000000000000000000000000;
                sprite[22] = 32'b00000000000000000000000000000000;
                sprite[23] = 32'b00000000000000000000000000000000;
                sprite[24] = 32'b00000000000000000000000000000000;
                sprite[25] = 32'b00000000000000000000000000000000;
                sprite[26] = 32'b00000000000000000000000000000000;
                sprite[27] = 32'b00000000000000000000000000000000;
                sprite[28] = 32'b00000000000000000000000000000000;
                sprite[29] = 32'b00000000000000000000000000000000;
                sprite[30] = 32'b00000000000000000000000000000000;
                sprite[31] = 32'b00000000000000000000000000000000;
				end
					 4'd5: begin
                sprite[0]  = 32'b00000000000000000000000000000000;
                sprite[1]  = 32'b00000000000000000000000000000000;
                sprite[2]  = 32'b00000000000000000000000000000000;
                sprite[3]  = 32'b00000000000000000000000000000000;
                sprite[4]  = 32'b00000000000000000000000000000000;
                sprite[5]  = 32'b00000000000000000000000000000000;
                sprite[6]  = 32'b00000000000000000000000000000000;
                sprite[7]  = 32'b00000000000000000000000000000000;
                sprite[8]  = 32'b00000000000000000000000000000000;
                sprite[9]  = 32'b00000000000000000000000000000000;
                sprite[10] = 32'b00000000000000000000000000000000;
                sprite[11] = 32'b00000000000000000000000000000000;
                sprite[12] = 32'b00000000000000000000000000000000;
                sprite[13] = 32'b00000000000000000000000000000000;
                sprite[14] = 32'b00000000000000000000000000000000;
                sprite[15] = 32'b00000000000000000000111110000000;
                sprite[16] = 32'b00000000000000000001111111000000;
                sprite[17] = 32'b00000000000000000111111111000000;
                sprite[18] = 32'b00000000000000000111111111000000;
                sprite[19] = 32'b00000000000000111111111111111000;
                sprite[20] = 32'b00000000000000111111111111111000;
                sprite[21] = 32'b00000000000011111111111111110000;
                sprite[22] = 32'b00000000000011111111111111110000;
                sprite[23] = 32'b00000000000111111111111111100000;
                sprite[24] = 32'b00000000000011111111111011000000;
                sprite[25] = 32'b00000000001111111111000000000000;
                sprite[26] = 32'b00000000001111000000000000000000;
                sprite[27] = 32'b00000000000000000000000000000000;
                sprite[28] = 32'b00000000000000000000000000000000;
                sprite[29] = 32'b00000000000000000000000000000000;
                sprite[30] = 32'b00000000000000000000000000000000;
                sprite[31] = 32'b00000000000000000000000000000000;
				end
					 4'd6: begin
                sprite[0]  = 32'b00000000000000000000000000000000;
                sprite[1]  = 32'b00000000000000000000000000000000;
                sprite[2]  = 32'b00000000000000000000000000000000;
                sprite[3]  = 32'b00000000000000000000000000000000;
                sprite[4]  = 32'b00000000000000000000000000000000;
                sprite[5]  = 32'b00000000000000000000000000000000;
                sprite[6]  = 32'b00000000000000000000000000000000;
                sprite[7]  = 32'b00000000000000000000000000000000;
                sprite[8]  = 32'b00000000000000000000000000000000;
                sprite[9]  = 32'b00000000000000000000000000000000;
                sprite[10] = 32'b00000000000000000000000000000000;
                sprite[11] = 32'b00000000000000000000000000000000;
                sprite[12] = 32'b00000000000000000000000000000000;
                sprite[13] = 32'b00000000000000000000000000000000;
                sprite[14] = 32'b00000000000000000000000000000000;
                sprite[15] = 32'b00000000000000000000001100000000;
                sprite[16] = 32'b00000000000000000000011110000000;
                sprite[17] = 32'b00000000000000000000111111000000;
                sprite[18] = 32'b00000000000000000000111111100000;
                sprite[19] = 32'b00000000000000000001111111110000;
                sprite[20] = 32'b00000000000000000011111111111000;
                sprite[21] = 32'b00000000000000000001111111111100;
                sprite[22] = 32'b00000000000000000011111111111100;
                sprite[23] = 32'b00000000000000000111111111111100;
                sprite[24] = 32'b00000000000000001111111111111000;
                sprite[25] = 32'b00000000000000001111111111010000;
                sprite[26] = 32'b00000000000000011111111110000000;
                sprite[27] = 32'b00000000000000011111111000000000;
                sprite[28] = 32'b00000000000000011110000000000000;
                sprite[29] = 32'b00000000000000001000000000000000;
                sprite[30] = 32'b00000000000000000000000000000000;
                sprite[31] = 32'b00000000000000000000000000000000;
				end
				

					 4'd7: begin
                sprite[0]  = 32'b00000000000000000000000000000000;
                sprite[1]  = 32'b00000000000000000000000000000000;
                sprite[2]  = 32'b00000000000000000000000000000000;
                sprite[3]  = 32'b00000000000000000000000000000000;
                sprite[4]  = 32'b00000000000000000000000000000000;
                sprite[5]  = 32'b00000000000000000000000000000000;
                sprite[6]  = 32'b00000000000000000000000000000000;
                sprite[7]  = 32'b00000000000000000000000000000000;
                sprite[8]  = 32'b00000000000000000000000000000000;
                sprite[9]  = 32'b00000000000000000000000000000000;
                sprite[10] = 32'b00000000000000000000000000000000;
                sprite[11] = 32'b00000000000001111000000000000000;
                sprite[12] = 32'b00000000000001111110000000000000;
                sprite[13] = 32'b00000000000011111111110000000000;
                sprite[14] = 32'b00000000000011111111111000000000;
                sprite[15] = 32'b00000000000001111111111000000000;
                sprite[16] = 32'b00000000000011111111111000000000;
                sprite[17] = 32'b00000000000011111111111000000000;
                sprite[18] = 32'b00000000000011111111110000000000;
                sprite[19] = 32'b00000000000011111111000000000000;
                sprite[20] = 32'b00000000000111111110000000000000;
                sprite[21] = 32'b00000000000011111100000000000000;
                sprite[22] = 32'b00000000000111111100000000000000;
                sprite[23] = 32'b00000000000111110100000000000000;
                sprite[24] = 32'b00000000000011110000000000000000;
                sprite[25] = 32'b00000000000111110000000000000000;
                sprite[26] = 32'b00000000000110000000000000000000;
                sprite[27] = 32'b00000000000000000000000000000000;
                sprite[28] = 32'b00000000000000000000000000000000;
                sprite[29] = 32'b00000000000000000000000000000000;
                sprite[30] = 32'b00000000000000000000000000000000;
                sprite[31] = 32'b00000000000000000000000000000000;
				end
					 4'd8: begin
                sprite[0]  = 32'b00000000000000000000000000000000;
                sprite[1]  = 32'b00000000000000000000000000000000;
                sprite[2]  = 32'b00000000000000000000000000000000;
                sprite[3]  = 32'b00000000000000000000000000000000;
                sprite[4]  = 32'b00000000000000000000000000000000;
                sprite[5]  = 32'b00000000000000000000000000000000;
                sprite[6]  = 32'b00000000000000000000000000000000;
                sprite[7]  = 32'b00000000000000000000000000000000;
                sprite[8]  = 32'b00000000000000000000000000000000;
                sprite[9]  = 32'b00000000000000000000000000000000;
                sprite[10] = 32'b00000000000111111111000000000000;
                sprite[11] = 32'b00000000001111111111100000000000;
                sprite[12] = 32'b00000000001111111111100000000000;
                sprite[13] = 32'b00000000001111111111100000000000;
                sprite[14] = 32'b00000000001111111111100000000000;
                sprite[15] = 32'b00000000000111111111000000000000;
                sprite[16] = 32'b00000000000111111111000000000000;
                sprite[17] = 32'b00000000000111111111000000000000;
                sprite[18] = 32'b00000000000011111110000000000000;
                sprite[19] = 32'b00000000000011111110000000000000;
                sprite[20] = 32'b00000000000011111110000000000000;
                sprite[21] = 32'b00000000000011111110000000000000;
                sprite[22] = 32'b00000000000001111100000000000000;
                sprite[23] = 32'b00000000000001111100000000000000;
                sprite[24] = 32'b00000000000001111100000000000000;
                sprite[25] = 32'b00000000000000111000000000000000;
                sprite[26] = 32'b00000000000000000000000000000000;
                sprite[27] = 32'b00000000000000000000000000000000;
                sprite[28] = 32'b00000000000000000000000000000000;
                sprite[29] = 32'b00000000000000000000000000000000;
                sprite[30] = 32'b00000000000000000000000000000000;
                sprite[31] = 32'b00000000000000000000000000000000;
				end
					 4'd9: begin
                sprite[0]  = 32'b00000000000000000000000000000000;
                sprite[1]  = 32'b00000000000000000000000000000000;
                sprite[2]  = 32'b00000000000000000000000000000000;
                sprite[3]  = 32'b00000000000000000000000000000000;
                sprite[4]  = 32'b00000000000000000000000000000000;
                sprite[5]  = 32'b00000000000000000000000000000000;
                sprite[6]  = 32'b00000000000000000000000000000000;
                sprite[7]  = 32'b00000000000000000000000000000000;
                sprite[8]  = 32'b00000000000000000000000000000000;
                sprite[9]  = 32'b00000000000000000000000000000000;
                sprite[10] = 32'b00000000000000000110000000000000;
                sprite[11] = 32'b00000000000000011111000000000000;
                sprite[12] = 32'b00000000000011111111100000000000;
                sprite[13] = 32'b00000000001111111111100000000000;
                sprite[14] = 32'b00000000001111111111000000000000;
                sprite[15] = 32'b00000000001111111111100000000000;
                sprite[16] = 32'b00000000001111111111100000000000;
                sprite[17] = 32'b00000000000111111111100000000000;
                sprite[18] = 32'b00000000000011111111100000000000;
                sprite[19] = 32'b00000000000001111111100000000000;
                sprite[20] = 32'b00000000000001111111110000000000;
                sprite[21] = 32'b00000000000000011111110000000000;
                sprite[22] = 32'b00000000000000011111100000000000;
                sprite[23] = 32'b00000000000000011111110000000000;
                sprite[24] = 32'b00000000000000000111110000000000;
                sprite[25] = 32'b00000000000000000011110000000000;
                sprite[26] = 32'b00000000000000000001100000000000;
                sprite[27] = 32'b00000000000000000000000000000000;
                sprite[28] = 32'b00000000000000000000000000000000;
                sprite[29] = 32'b00000000000000000000000000000000;
                sprite[30] = 32'b00000000000000000000000000000000;
                sprite[31] = 32'b00000000000000000000000000000000;
				end
            4'd10: begin
                sprite[0]  = 32'b00000000000000000000000000000000;
                sprite[1]  = 32'b00000000000000000000000000000000;
                sprite[2]  = 32'b00000000000000000000000000000000;
                sprite[3]  = 32'b00000000000000000000000000000000;
                sprite[4]  = 32'b00000000000000000000000000000000;
                sprite[5]  = 32'b00000000000000000000000000000000;
                sprite[6]  = 32'b00000000000000000000000000000000;
                sprite[7]  = 32'b00000000000000000000000000000000;
                sprite[8]  = 32'b00000000000000000000000000000000;
                sprite[9]  = 32'b00000000000000000000000000000000;
                sprite[10] = 32'b00000000000000000000000000000000;
                sprite[11] = 32'b00000000000000000000000000000000;
                sprite[12] = 32'b00000000000000000111000000000000;
                sprite[13] = 32'b00000000000000001111100000000000;
                sprite[14] = 32'b00000000000000011111110000000000;
                sprite[15] = 32'b00000000000000111111100000000000;
                sprite[16] = 32'b00000000000001111111110000000000;
                sprite[17] = 32'b00000000000011111111111000000000;
                sprite[18] = 32'b00000000000111111111111000000000;
                sprite[19] = 32'b00000000000111111111111100000000;
                sprite[20] = 32'b00000000000011111111111110000000;
                sprite[21] = 32'b00000000000001111111111110000000;
                sprite[22] = 32'b00000000000000011111111110000000;
                sprite[23] = 32'b00000000000000001111111111000000;
                sprite[24] = 32'b00000000000000000001111111000000;
                sprite[25] = 32'b00000000000000000000111111100000;
                sprite[26] = 32'b00000000000000000000001111000000;
                sprite[27] = 32'b00000000000000000000000000000000;
                sprite[28] = 32'b00000000000000000000000000000000;
                sprite[29] = 32'b00000000000000000000000000000000;
                sprite[30] = 32'b00000000000000000000000000000000;
                sprite[31] = 32'b00000000000000000000000000000000;
            end
            4'd11: begin
                sprite[0]  = 32'b00000000000000000000000000000000;
                sprite[1]  = 32'b00000000000000000000000000000000;
                sprite[2]  = 32'b00000000000000000000000000000000;
                sprite[3]  = 32'b00000000000000000000000000000000;
                sprite[4]  = 32'b00000000000000000000000000000000;
                sprite[5]  = 32'b00000000000000000000000000000000;
                sprite[6]  = 32'b00000000000000000000000000000000;
                sprite[7]  = 32'b00000000000000000000000000000000;
                sprite[8]  = 32'b00000000000000000000000000000000;
                sprite[9]  = 32'b00000000000000000000000000000000;
                sprite[10] = 32'b00000000000000000000000000000000;
                sprite[11] = 32'b00000000000001111000000000000000;
                sprite[12] = 32'b00000000000011111100000000000000;
                sprite[13] = 32'b00000000000011111110000000000000;
                sprite[14] = 32'b00000000000011111111000000000000;
                sprite[15] = 32'b00000000000111111111100000000000;
                sprite[16] = 32'b00000000000111111111111100000000;
                sprite[17] = 32'b00000000001111111111111000000000;
                sprite[18] = 32'b00000000001111111111111111000000;
                sprite[19] = 32'b00000000001111111111111111000000;
                sprite[20] = 32'b00000000001111111111111111000000;
                sprite[21] = 32'b00000000000011011111111111000000;
                sprite[22] = 32'b00000000000000000000101101100000;
                sprite[23] = 32'b00000000000000000000000001100000;
                sprite[24] = 32'b00000000000000000000000000000000;
                sprite[25] = 32'b00000000000000000000000000000000;
                sprite[26] = 32'b00000000000000000000000000000000;
                sprite[27] = 32'b00000000000000000000000000000000;
                sprite[28] = 32'b00000000000000000000000000000000;
                sprite[29] = 32'b00000000000000000000000000000000;
                sprite[30] = 32'b00000000000000000000000000000000;
                sprite[31] = 32'b00000000000000000000000000000000;
            end
            4'd12: begin
                sprite[0]  = 32'b00000000000000000000000000000000;
                sprite[1]  = 32'b00000000000000000000000000000000;
                sprite[2]  = 32'b00000000000000000000000000000000;
                sprite[3]  = 32'b00000000000000000000000000000000;
                sprite[4]  = 32'b00000000000000000000000000000000;
                sprite[5]  = 32'b00000000000000000000000000000000;
                sprite[6]  = 32'b00000000000000000000000000000000;
                sprite[7]  = 32'b00000000000000000000000000000000;
                sprite[8]  = 32'b00000000000000000000000000000000;
                sprite[9]  = 32'b00000000000000000000000000000000;
                sprite[10] = 32'b00000000000000000000000000000000;
                sprite[11] = 32'b00000000000111100000000000000000;
                sprite[12] = 32'b00000000001111111100000000000000;
                sprite[13] = 32'b00000000001111111111110000000000;
                sprite[14] = 32'b00000000001111111111111111000000;
                sprite[15] = 32'b00000000001111111111111111000000;
                sprite[16] = 32'b00000000001111111111111111000000;
                sprite[17] = 32'b00000000001111111111111110000000;
                sprite[18] = 32'b00000000001111111111110000000000;
                sprite[19] = 32'b00000000001111111100000000000000;
                sprite[20] = 32'b00000000000111100000000000000000;
                sprite[21] = 32'b00000000000000000000000000000000;
                sprite[22] = 32'b00000000000000000000000000000000;
                sprite[23] = 32'b00000000000000000000000000000000;
                sprite[24] = 32'b00000000000000000000000000000000;
                sprite[25] = 32'b00000000000000000000000000000000;
                sprite[26] = 32'b00000000000000000000000000000000;
                sprite[27] = 32'b00000000000000000000000000000000;
                sprite[28] = 32'b00000000000000000000000000000000;
                sprite[29] = 32'b00000000000000000000000000000000;
                sprite[30] = 32'b00000000000000000000000000000000;
                sprite[31] = 32'b00000000000000000000000000000000;
            end
            4'd13: begin
                sprite[0]  = 32'b00000000000000000000000000000000;
                sprite[1]  = 32'b00000000000000000000000000000000;
                sprite[2]  = 32'b00000000000000000000000000000000;
                sprite[3]  = 32'b00000000000000000000000000000000;
                sprite[4]  = 32'b00000000000000000000000000000000;
                sprite[5]  = 32'b00000000000000000000000000000000;
                sprite[6]  = 32'b00000000000000000000000000000000;
                sprite[7]  = 32'b00000000000000000000000000000000;
                sprite[8]  = 32'b00000000000000000000000000000000;
                sprite[9]  = 32'b00000000000000000000000001100000;
                sprite[10] = 32'b00000000000000000000110111100000;
                sprite[11] = 32'b00000000000011011111111111000000;
                sprite[12] = 32'b00000000000111111111111111100000;
                sprite[13] = 32'b00000000001111111111111111000000;
                sprite[14] = 32'b00000000001111111111111111000000;
                sprite[15] = 32'b00000000000111111111111100000000;
                sprite[16] = 32'b00000000000111111111111100000000;
                sprite[17] = 32'b00000000000011111111100000000000;
                sprite[18] = 32'b00000000000011111111100000000000;
                sprite[19] = 32'b00000000000011111110000000000000;
                sprite[20] = 32'b00000000000001111100000000000000;
                sprite[21] = 32'b00000000000001111000000000000000;
                sprite[22] = 32'b00000000000000000000000000000000;
                sprite[23] = 32'b00000000000000000000000000000000;
                sprite[24] = 32'b00000000000000000000000000000000;
                sprite[25] = 32'b00000000000000000000000000000000;
                sprite[26] = 32'b00000000000000000000000000000000;
                sprite[27] = 32'b00000000000000000000000000000000;
                sprite[28] = 32'b00000000000000000000000000000000;
                sprite[29] = 32'b00000000000000000000000000000000;
                sprite[30] = 32'b00000000000000000000000000000000;
                sprite[31] = 32'b00000000000000000000000000000000;
            end
            4'd14: begin
                sprite[0]  = 32'b00000000000000000000000000000000;
                sprite[1]  = 32'b00000000000000000000000000000000;
                sprite[2]  = 32'b00000000000000000000000000000000;
                sprite[3]  = 32'b00000000000000000000000000000000;
                sprite[4]  = 32'b00000000000000000000000000000000;
                sprite[5]  = 32'b00000000000000000000000000000000;
                sprite[6]  = 32'b00000000000000000000000000000000;
                sprite[7]  = 32'b00000000000000000000000000000000;
                sprite[8]  = 32'b00000000000000000000000000000000;
                sprite[9]  = 32'b00000000000000000000000001000000;
                sprite[10] = 32'b00000000000000000000000111100000;
                sprite[11] = 32'b00000000000000000000111111100000;
                sprite[12] = 32'b00000000000000000001111111100000;
                sprite[13] = 32'b00000000000000000111111111100000;
                sprite[14] = 32'b00000000000000101111111111000000;
                sprite[15] = 32'b00000000000001111111111111000000;
                sprite[16] = 32'b00000000000011111111111110000000;
                sprite[17] = 32'b00000000000011111111111100000000;
                sprite[18] = 32'b00000000000011111111111000000000;
                sprite[19] = 32'b00000000000001111111111100000000;
                sprite[20] = 32'b00000000000000111111111000000000;
                sprite[21] = 32'b00000000000000011111110000000000;
                sprite[22] = 32'b00000000000000001111110000000000;
                sprite[23] = 32'b00000000000000000111100000000000;
                sprite[24] = 32'b00000000000000000011000000000000;
                sprite[25] = 32'b00000000000000000000000000000000;
                sprite[26] = 32'b00000000000000000000000000000000;
                sprite[27] = 32'b00000000000000000000000000000000;
                sprite[28] = 32'b00000000000000000000000000000000;
                sprite[29] = 32'b00000000000000000000000000000000;
                sprite[30] = 32'b00000000000000000000000000000000;
                sprite[31] = 32'b00000000000000000000000000000000;
            end
            4'd15: begin
                sprite[0]  = 32'b00000000000000000000000000000000;
                sprite[1]  = 32'b00000000000000000000000000000000;
                sprite[2]  = 32'b00000000000000000000000000000000;
                sprite[3]  = 32'b00000000000000000000000000000000;
                sprite[4]  = 32'b00000000000000000000000000000000;
                sprite[5]  = 32'b00000000000000000000000000000000;
                sprite[6]  = 32'b00000000000000000000000000000000;
                sprite[7]  = 32'b00000000000000000000000000000000;
                sprite[8]  = 32'b00000000000000000001111000000000;
                sprite[9]  = 32'b00000000000000000011111000000000;
                sprite[10] = 32'b00000000000000000111111000000000;
                sprite[11] = 32'b00000000000000001111111000000000;
                sprite[12] = 32'b00000000000000001111110000000000;
                sprite[13] = 32'b00000000000000011111111000000000;
                sprite[14] = 32'b00000000000000111111110000000000;
                sprite[15] = 32'b00000000000001111111110000000000;
                sprite[16] = 32'b00000000000011111111110000000000;
                sprite[17] = 32'b00000000000111111111110000000000;
                sprite[18] = 32'b00000000001111111111110000000000;
                sprite[19] = 32'b00000000001111111111100000000000;
                sprite[20] = 32'b00000000001111111111110000000000;
                sprite[21] = 32'b00000000011111111111110000000000;
                sprite[22] = 32'b00000000000000111111100000000000;
                sprite[23] = 32'b00000000000000001111100000000000;
                sprite[24] = 32'b00000000000000000000000000000000;
                sprite[25] = 32'b00000000000000000000000000000000;
                sprite[26] = 32'b00000000000000000000000000000000;
                sprite[27] = 32'b00000000000000000000000000000000;
                sprite[28] = 32'b00000000000000000000000000000000;
                sprite[29] = 32'b00000000000000000000000000000000;
                sprite[30] = 32'b00000000000000000000000000000000;
                sprite[31] = 32'b00000000000000000000000000000000;
            end				
			endcase
	end
    wire signed [9:0] x_rel, y_rel;
    assign x_rel = hcount - x_center;
    assign y_rel = vcount - y_center;

    always @(*) begin
        // Default color is black
        rgb = 24'h000000;
        // Check if the current pixel is within the bounds of the sprite
        if (x_rel >= -16 && x_rel < 16 && y_rel >= -16 && y_rel < 16) begin
            if (sprite[y_rel + 16][x_rel + 16]) begin
                rgb = 24'hFFFFFF; // White color for the player sprite
            end
        end
    end
endmodule


