module shooting_name(
input [9:0] hsync,
input [9:0] vsync,
output reg [23:0] rgb );

reg [0:159] sprite [0:39];

always @(*) begin


sprite[0] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[1] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[2] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[3] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[4] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[5] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[6] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[7] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[8] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[9] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[10] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[11] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[12] =  160'b0000000000000000000000011000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[13] =  160'b0001111110000000000000011000000000000000000000000000000000000000000000011000000011000001110000001100000000000000000000000000000000000000000000000000000000000000;
sprite[14] =  160'b0011100110000000000000011000000000000000000000001000000000000000000000011000000011000001110000011000000000000000000000000000000000000000000000000000000000000000;
sprite[15] =  160'b0011000000000000000000011000000000000000000000001000000000000000000000011000000011000001110000011000000000000000000000000000000000000000000000000000000000000000;
sprite[16] =  160'b0011000000000011110000011000001110000000111100111111000011110000000111011000000001100001011000011000011110000001111000001001110000000111100000110111100000110000;
sprite[17] =  160'b0011000000000111111000011000111111100001111110111111000111111000011111111000000001100011011000010000111111000011111100001011111000001111111000111111110000110000;
sprite[18] =  160'b0001110000001100001100011000100001100011000010001000001100001100011000111000000001100011011000110001100001100100000110001100001100011000011000111000110000110000;
sprite[19] =  160'b0000111100001000001100011001100000110011000000001000001100000100110000011000000000100011001000110001000001100000000110001100001100011000001100110000010000000000;
sprite[20] =  160'b0000001110011111111100011001111111110011000000001000001111111100110000011000000000110010001100110011111111100000111110001100001100110000001100110000010000000000;
sprite[21] =  160'b0000000011011111111100011001111111100011000000001000001111111100110000011000000000110110001101100011111111100011111110001100000100110000001100110000010000000000;
sprite[22] =  160'b0000000011011000000000011001100000000011000000001000001100000000110000011000000000110110001101100011000000000110000110001100001100110000001100110000010000000000;
sprite[23] =  160'b0000000011001100000000011001100000000011000000001000001100000000111000011000000000011110000111100001100000000110000110001100001100011000001100110000010000000000;
sprite[24] =  160'b0111001110001110000100011000110000100011100110001101000110000100011001111000000000011100000111000001110000100110001110001110011100011100111000110000010000110000;
sprite[25] =  160'b0011111100000111111100011000011111100001111110001111000111111100001111011000000000011100000111000000111111100011111110001111111000001111110000110000010000110000;
sprite[26] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000;
sprite[27] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000;
sprite[28] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000;
sprite[29] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000;
sprite[30] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[31] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[32] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[33] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[34] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[35] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[36] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[37] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[38] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
sprite[39] =  160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

end




wire signed [9:0] x_rel, y_rel;
assign x_rel = hsync - 560;
assign y_rel = vsync - 390;

    always @(*) begin
        if (x_rel >= -80 && x_rel < 80 && y_rel >= -20 && y_rel < 20) begin
            if (sprite[y_rel + 20][x_rel + 80]) begin
                rgb = 24'hFFFF00;
				end
				else begin 
				rgb = 24'h000000;
				end
			end
			else begin
			rgb =24'h000000;
		end
    end
endmodule

