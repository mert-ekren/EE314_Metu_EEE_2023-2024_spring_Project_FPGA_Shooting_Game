module yzler(
input [3:0] digit100,
input [9:0] hsync,
input [9:0] vsync,
output reg [23:0] rgb
);

reg [0:49] sprite [0:49];

always @(*) begin

	case (digit100) 
		4'd0: begin
sprite[0] =  50'b00000000000000000000000000000000000000000000000000;
sprite[1] =  50'b00000000000000000000000000000000000000000000000000;
sprite[2] =  50'b00000000000000000000000000000000000000000000000000;
sprite[3] =  50'b00000000000000000000000000000000000000000000000000;
sprite[4] =  50'b00000000000000000000000000000000000000000000000000;
sprite[5] =  50'b00000000000000000000000000000000000000000000000000;
sprite[6] =  50'b00000000000000000000000000000000000000000000000000;
sprite[7] =  50'b00000000000000000000000000000000000000000000000000;
sprite[8] =  50'b00000000000000000000000000000000000000000000000000;
sprite[9] =  50'b00000000000000000000000000000000000000000000000000;
sprite[10] =  50'b00000000000000000000000000000000000000000000000000;
sprite[11] =  50'b00000000000000000000000000000000000000000000000000;
sprite[12] =  50'b00000000000000000000000000000000000000000000000000;
sprite[13] =  50'b00000000000000000000000000000000000000000000000000;
sprite[14] =  50'b00000000000000000000000110000000000000000000000000;
sprite[15] =  50'b00000000000000000000111111110000000000000000000000;
sprite[16] =  50'b00000000000000000001111111111000000000000000000000;
sprite[17] =  50'b00000000000000000011110000111100000000000000000000;
sprite[18] =  50'b00000000000000000111100000011100000000000000000000;
sprite[19] =  50'b00000000000000000111000000011110000000000000000000;
sprite[20] =  50'b00000000000000000111000000001110000000000000000000;
sprite[21] =  50'b00000000000000001111000000001110000000000000000000;
sprite[22] =  50'b00000000000000001110000000001110000000000000000000;
sprite[23] =  50'b00000000000000001110000000001110000000000000000000;
sprite[24] =  50'b00000000000000001110000000001110000000000000000000;
sprite[25] =  50'b00000000000000001110000000001110000000000000000000;
sprite[26] =  50'b00000000000000001110000000001110000000000000000000;
sprite[27] =  50'b00000000000000001110000000001110000000000000000000;
sprite[28] =  50'b00000000000000001110000000001110000000000000000000;
sprite[29] =  50'b00000000000000001110000000001110000000000000000000;
sprite[30] =  50'b00000000000000001111000000001110000000000000000000;
sprite[31] =  50'b00000000000000000111000000001110000000000000000000;
sprite[32] =  50'b00000000000000000111000000011110000000000000000000;
sprite[33] =  50'b00000000000000000111100000011100000000000000000000;
sprite[34] =  50'b00000000000000000011110000111100000000000000000000;
sprite[35] =  50'b00000000000000000011111111111000000000000000000000;
sprite[36] =  50'b00000000000000000000111111110000000000000000000000;
sprite[37] =  50'b00000000000000000000001110000000000000000000000000;
sprite[38] =  50'b00000000000000000000000000000000000000000000000000;
sprite[39] =  50'b00000000000000000000000000000000000000000000000000;
sprite[40] =  50'b00000000000000000000000000000000000000000000000000;
sprite[41] =  50'b00000000000000000000000000000000000000000000000000;
sprite[42] =  50'b00000000000000000000000000000000000000000000000000;
sprite[43] =  50'b00000000000000000000000000000000000000000000000000;
sprite[44] =  50'b00000000000000000000000000000000000000000000000000;
sprite[45] =  50'b00000000000000000000000000000000000000000000000000;
sprite[46] =  50'b00000000000000000000000000000000000000000000000000;
sprite[47] =  50'b00000000000000000000000000000000000000000000000000;
sprite[48] =  50'b00000000000000000000000000000000000000000000000000;
sprite[49] =  50'b00000000000000000000000000000000000000000000000000;
		end
		
		4'd1: begin
sprite[0] =  50'b00000000000000000000000000000000000000000000000000;
sprite[1] =  50'b00000000000000000000000000000000000000000000000000;
sprite[2] =  50'b00000000000000000000000000000000000000000000000000;
sprite[3] =  50'b00000000000000000000000000000000000000000000000000;
sprite[4] =  50'b00000000000000000000000000000000000000000000000000;
sprite[5] =  50'b00000000000000000000000000000000000000000000000000;
sprite[6] =  50'b00000000000000000000000000000000000000000000000000;
sprite[7] =  50'b00000000000000000000000000000000000000000000000000;
sprite[8] =  50'b00000000000000000000000000000000000000000000000000;
sprite[9] =  50'b00000000000000000000000000000000000000000000000000;
sprite[10] =  50'b00000000000000000000000000000000000000000000000000;
sprite[11] =  50'b00000000000000000000000000000000000000000000000000;
sprite[12] =  50'b00000000000000000000000000000000000000000000000000;
sprite[13] =  50'b00000000000000000000000000000000000000000000000000;
sprite[14] =  50'b00000000000000000000000000000000000000000000000000;
sprite[15] =  50'b00000000000000000000000111000000000000000000000000;
sprite[16] =  50'b00000000000000000000011111000000000000000000000000;
sprite[17] =  50'b00000000000000000000111111000000000000000000000000;
sprite[18] =  50'b00000000000000000011111111000000000000000000000000;
sprite[19] =  50'b00000000000000000011100111000000000000000000000000;
sprite[20] =  50'b00000000000000000010000111000000000000000000000000;
sprite[21] =  50'b00000000000000000000000111000000000000000000000000;
sprite[22] =  50'b00000000000000000000000111000000000000000000000000;
sprite[23] =  50'b00000000000000000000000111000000000000000000000000;
sprite[24] =  50'b00000000000000000000000111000000000000000000000000;
sprite[25] =  50'b00000000000000000000000111000000000000000000000000;
sprite[26] =  50'b00000000000000000000000111000000000000000000000000;
sprite[27] =  50'b00000000000000000000000111000000000000000000000000;
sprite[28] =  50'b00000000000000000000000111000000000000000000000000;
sprite[29] =  50'b00000000000000000000000111000000000000000000000000;
sprite[30] =  50'b00000000000000000000000111000000000000000000000000;
sprite[31] =  50'b00000000000000000000000111000000000000000000000000;
sprite[32] =  50'b00000000000000000000000111000000000000000000000000;
sprite[33] =  50'b00000000000000000000000111000000000000000000000000;
sprite[34] =  50'b00000000000000000000001111000000000000000000000000;
sprite[35] =  50'b00000000000000000011111111111110000000000000000000;
sprite[36] =  50'b00000000000000000011111111111110000000000000000000;
sprite[37] =  50'b00000000000000000000000000000000000000000000000000;
sprite[38] =  50'b00000000000000000000000000000000000000000000000000;
sprite[39] =  50'b00000000000000000000000000000000000000000000000000;
sprite[40] =  50'b00000000000000000000000000000000000000000000000000;
sprite[41] =  50'b00000000000000000000000000000000000000000000000000;
sprite[42] =  50'b00000000000000000000000000000000000000000000000000;
sprite[43] =  50'b00000000000000000000000000000000000000000000000000;
sprite[44] =  50'b00000000000000000000000000000000000000000000000000;
sprite[45] =  50'b00000000000000000000000000000000000000000000000000;
sprite[46] =  50'b00000000000000000000000000000000000000000000000000;
sprite[47] =  50'b00000000000000000000000000000000000000000000000000;
sprite[48] =  50'b00000000000000000000000000000000000000000000000000;
sprite[49] =  50'b00000000000000000000000000000000000000000000000000;
		end
		
		4'd2: begin
sprite[0] =  50'b00000000000000000000000000000000000000000000000000;
sprite[1] =  50'b00000000000000000000000000000000000000000000000000;
sprite[2] =  50'b00000000000000000000000000000000000000000000000000;
sprite[3] =  50'b00000000000000000000000000000000000000000000000000;
sprite[4] =  50'b00000000000000000000000000000000000000000000000000;
sprite[5] =  50'b00000000000000000000000000000000000000000000000000;
sprite[6] =  50'b00000000000000000000000000000000000000000000000000;
sprite[7] =  50'b00000000000000000000000000000000000000000000000000;
sprite[8] =  50'b00000000000000000000000000000000000000000000000000;
sprite[9] =  50'b00000000000000000000000000000000000000000000000000;
sprite[10] =  50'b00000000000000000000000000000000000000000000000000;
sprite[11] =  50'b00000000000000000000000000000000000000000000000000;
sprite[12] =  50'b00000000000000000000000000000000000000000000000000;
sprite[13] =  50'b00000000000000000000000000000000000000000000000000;
sprite[14] =  50'b00000000000000000000000110000000000000000000000000;
sprite[15] =  50'b00000000000000000000111111110000000000000000000000;
sprite[16] =  50'b00000000000000000011111111111000000000000000000000;
sprite[17] =  50'b00000000000000000011110001111100000000000000000000;
sprite[18] =  50'b00000000000000000011000000111100000000000000000000;
sprite[19] =  50'b00000000000000000000000000011110000000000000000000;
sprite[20] =  50'b00000000000000000000000000011110000000000000000000;
sprite[21] =  50'b00000000000000000000000000011100000000000000000000;
sprite[22] =  50'b00000000000000000000000000011100000000000000000000;
sprite[23] =  50'b00000000000000000000000000011100000000000000000000;
sprite[24] =  50'b00000000000000000000000000111100000000000000000000;
sprite[25] =  50'b00000000000000000000000000111000000000000000000000;
sprite[26] =  50'b00000000000000000000000001110000000000000000000000;
sprite[27] =  50'b00000000000000000000000011110000000000000000000000;
sprite[28] =  50'b00000000000000000000000111100000000000000000000000;
sprite[29] =  50'b00000000000000000000000111000000000000000000000000;
sprite[30] =  50'b00000000000000000000001110000000000000000000000000;
sprite[31] =  50'b00000000000000000000011100000000000000000000000000;
sprite[32] =  50'b00000000000000000000111000000000000000000000000000;
sprite[33] =  50'b00000000000000000001110000000000000000000000000000;
sprite[34] =  50'b00000000000000000011111111111110000000000000000000;
sprite[35] =  50'b00000000000000000011111111111110000000000000000000;
sprite[36] =  50'b00000000000000000011111111111110000000000000000000;
sprite[37] =  50'b00000000000000000000000000000000000000000000000000;
sprite[38] =  50'b00000000000000000000000000000000000000000000000000;
sprite[39] =  50'b00000000000000000000000000000000000000000000000000;
sprite[40] =  50'b00000000000000000000000000000000000000000000000000;
sprite[41] =  50'b00000000000000000000000000000000000000000000000000;
sprite[42] =  50'b00000000000000000000000000000000000000000000000000;
sprite[43] =  50'b00000000000000000000000000000000000000000000000000;
sprite[44] =  50'b00000000000000000000000000000000000000000000000000;
sprite[45] =  50'b00000000000000000000000000000000000000000000000000;
sprite[46] =  50'b00000000000000000000000000000000000000000000000000;
sprite[47] =  50'b00000000000000000000000000000000000000000000000000;
sprite[48] =  50'b00000000000000000000000000000000000000000000000000;
sprite[49] =  50'b00000000000000000000000000000000000000000000000000;

		end
		
		4'd3: begin
sprite[0] =  50'b00000000000000000000000000000000000000000000000000;
sprite[1] =  50'b00000000000000000000000000000000000000000000000000;
sprite[2] =  50'b00000000000000000000000000000000000000000000000000;
sprite[3] =  50'b00000000000000000000000000000000000000000000000000;
sprite[4] =  50'b00000000000000000000000000000000000000000000000000;
sprite[5] =  50'b00000000000000000000000000000000000000000000000000;
sprite[6] =  50'b00000000000000000000000000000000000000000000000000;
sprite[7] =  50'b00000000000000000000000000000000000000000000000000;
sprite[8] =  50'b00000000000000000000000000000000000000000000000000;
sprite[9] =  50'b00000000000000000000000000000000000000000000000000;
sprite[10] =  50'b00000000000000000000000000000000000000000000000000;
sprite[11] =  50'b00000000000000000000001100000000000000000000000000;
sprite[12] =  50'b00000000000000000001111111100000000000000000000000;
sprite[13] =  50'b00000000000000000011111111110000000000000000000000;
sprite[14] =  50'b00000000000000000111100001111000000000000000000000;
sprite[15] =  50'b00000000000000000110000000111000000000000000000000;
sprite[16] =  50'b00000000000000000000000000111000000000000000000000;
sprite[17] =  50'b00000000000000000000000000111000000000000000000000;
sprite[18] =  50'b00000000000000000000000000111000000000000000000000;
sprite[19] =  50'b00000000000000000000000000111000000000000000000000;
sprite[20] =  50'b00000000000000000000000001111000000000000000000000;
sprite[21] =  50'b00000000000000000000000111110000000000000000000000;
sprite[22] =  50'b00000000000000000001111111000000000000000000000000;
sprite[23] =  50'b00000000000000000001111111110000000000000000000000;
sprite[24] =  50'b00000000000000000000000011111000000000000000000000;
sprite[25] =  50'b00000000000000000000000000111100000000000000000000;
sprite[26] =  50'b00000000000000000000000000011100000000000000000000;
sprite[27] =  50'b00000000000000000000000000011100000000000000000000;
sprite[28] =  50'b00000000000000000000000000011100000000000000000000;
sprite[29] =  50'b00000000000000000000000000011100000000000000000000;
sprite[30] =  50'b00000000000000000000000000111100000000000000000000;
sprite[31] =  50'b00000000000000000111000001111000000000000000000000;
sprite[32] =  50'b00000000000000000111111111111000000000000000000000;
sprite[33] =  50'b00000000000000000011111111100000000000000000000000;
sprite[34] =  50'b00000000000000000000001100000000000000000000000000;
sprite[35] =  50'b00000000000000000000000000000000000000000000000000;
sprite[36] =  50'b00000000000000000000000000000000000000000000000000;
sprite[37] =  50'b00000000000000000000000000000000000000000000000000;
sprite[38] =  50'b00000000000000000000000000000000000000000000000000;
sprite[39] =  50'b00000000000000000000000000000000000000000000000000;
sprite[40] =  50'b00000000000000000000000000000000000000000000000000;
sprite[41] =  50'b00000000000000000000000000000000000000000000000000;
sprite[42] =  50'b00000000000000000000000000000000000000000000000000;
sprite[43] =  50'b00000000000000000000000000000000000000000000000000;
sprite[44] =  50'b00000000000000000000000000000000000000000000000000;
sprite[45] =  50'b00000000000000000000000000000000000000000000000000;
sprite[46] =  50'b00000000000000000000000000000000000000000000000000;
sprite[47] =  50'b00000000000000000000000000000000000000000000000000;
sprite[48] =  50'b00000000000000000000000000000000000000000000000000;
sprite[49] =  50'b00000000000000000000000000000000000000000000000000;
		
		end
		
		4'd4: begin
sprite[0] =  50'b00000000000000000000000000000000000000000000000000;
sprite[1] =  50'b00000000000000000000000000000000000000000000000000;
sprite[2] =  50'b00000000000000000000000000000000000000000000000000;
sprite[3] =  50'b00000000000000000000000000000000000000000000000000;
sprite[4] =  50'b00000000000000000000000000000000000000000000000000;
sprite[5] =  50'b00000000000000000000000000000000000000000000000000;
sprite[6] =  50'b00000000000000000000000000000000000000000000000000;
sprite[7] =  50'b00000000000000000000000000000000000000000000000000;
sprite[8] =  50'b00000000000000000000000000000000000000000000000000;
sprite[9] =  50'b00000000000000000000000000000000000000000000000000;
sprite[10] =  50'b00000000000000000000000000000000000000000000000000;
sprite[11] =  50'b00000000000000000000000000000000000000000000000000;
sprite[12] =  50'b00000000000000000000000000000000000000000000000000;
sprite[13] =  50'b00000000000000000000000000000000000000000000000000;
sprite[14] =  50'b00000000000000000000000001111000000000000000000000;
sprite[15] =  50'b00000000000000000000000011111000000000000000000000;
sprite[16] =  50'b00000000000000000000000011111000000000000000000000;
sprite[17] =  50'b00000000000000000000000111111000000000000000000000;
sprite[18] =  50'b00000000000000000000000110011000000000000000000000;
sprite[19] =  50'b00000000000000000000001110011000000000000000000000;
sprite[20] =  50'b00000000000000000000011100011000000000000000000000;
sprite[21] =  50'b00000000000000000000011100011000000000000000000000;
sprite[22] =  50'b00000000000000000000111000011000000000000000000000;
sprite[23] =  50'b00000000000000000000111000011000000000000000000000;
sprite[24] =  50'b00000000000000000001110000011000000000000000000000;
sprite[25] =  50'b00000000000000000001100000011000000000000000000000;
sprite[26] =  50'b00000000000000000011100000011000000000000000000000;
sprite[27] =  50'b00000000000000000111000000011000000000000000000000;
sprite[28] =  50'b00000000000000000111000000111100000000000000000000;
sprite[29] =  50'b00000000000000000111111111111111100000000000000000;
sprite[30] =  50'b00000000000000000111111111111111000000000000000000;
sprite[31] =  50'b00000000000000000000000000011000000000000000000000;
sprite[32] =  50'b00000000000000000000000000011000000000000000000000;
sprite[33] =  50'b00000000000000000000000000011000000000000000000000;
sprite[34] =  50'b00000000000000000000000000011000000000000000000000;
sprite[35] =  50'b00000000000000000000000000011000000000000000000000;
sprite[36] =  50'b00000000000000000000000000000000000000000000000000;
sprite[37] =  50'b00000000000000000000000000000000000000000000000000;
sprite[38] =  50'b00000000000000000000000000000000000000000000000000;
sprite[39] =  50'b00000000000000000000000000000000000000000000000000;
sprite[40] =  50'b00000000000000000000000000000000000000000000000000;
sprite[41] =  50'b00000000000000000000000000000000000000000000000000;
sprite[42] =  50'b00000000000000000000000000000000000000000000000000;
sprite[43] =  50'b00000000000000000000000000000000000000000000000000;
sprite[44] =  50'b00000000000000000000000000000000000000000000000000;
sprite[45] =  50'b00000000000000000000000000000000000000000000000000;
sprite[46] =  50'b00000000000000000000000000000000000000000000000000;
sprite[47] =  50'b00000000000000000000000000000000000000000000000000;
sprite[48] =  50'b00000000000000000000000000000000000000000000000000;
sprite[49] =  50'b00000000000000000000000000000000000000000000000000;
		
		end
		
		4'd5: begin
sprite[0] =  50'b00000000000000000000000000000000000000000000000000;
sprite[1] =  50'b00000000000000000000000000000000000000000000000000;
sprite[2] =  50'b00000000000000000000000000000000000000000000000000;
sprite[3] =  50'b00000000000000000000000000000000000000000000000000;
sprite[4] =  50'b00000000000000000000000000000000000000000000000000;
sprite[5] =  50'b00000000000000000000000000000000000000000000000000;
sprite[6] =  50'b00000000000000000000000000000000000000000000000000;
sprite[7] =  50'b00000000000000000000000000000000000000000000000000;
sprite[8] =  50'b00000000000000000000000000000000000000000000000000;
sprite[9] =  50'b00000000000000000000000000000000000000000000000000;
sprite[10] =  50'b00000000000000000000000000000000000000000000000000;
sprite[11] =  50'b00000000000000000000000000000000000000000000000000;
sprite[12] =  50'b00000000000000000000000000000000000000000000000000;
sprite[13] =  50'b00000000000000000000000000000000000000000000000000;
sprite[14] =  50'b00000000000000000000000000000000000000000000000000;
sprite[15] =  50'b00000000000000000000111111111110000000000000000000;
sprite[16] =  50'b00000000000000000000111111111110000000000000000000;
sprite[17] =  50'b00000000000000000000111111111100000000000000000000;
sprite[18] =  50'b00000000000000000000110000000000000000000000000000;
sprite[19] =  50'b00000000000000000000110000000000000000000000000000;
sprite[20] =  50'b00000000000000000000110000000000000000000000000000;
sprite[21] =  50'b00000000000000000000110000000000000000000000000000;
sprite[22] =  50'b00000000000000000000110000000000000000000000000000;
sprite[23] =  50'b00000000000000000000111000000000000000000000000000;
sprite[24] =  50'b00000000000000000000111111111000000000000000000000;
sprite[25] =  50'b00000000000000000000111111111110000000000000000000;
sprite[26] =  50'b00000000000000000000000000011110000000000000000000;
sprite[27] =  50'b00000000000000000000000000001111000000000000000000;
sprite[28] =  50'b00000000000000000000000000000111000000000000000000;
sprite[29] =  50'b00000000000000000000000000000111100000000000000000;
sprite[30] =  50'b00000000000000000000000000000111100000000000000000;
sprite[31] =  50'b00000000000000000000000000000111000000000000000000;
sprite[32] =  50'b00000000000000000000000000000111000000000000000000;
sprite[33] =  50'b00000000000000000000000000001111000000000000000000;
sprite[34] =  50'b00000000000000000001100000011110000000000000000000;
sprite[35] =  50'b00000000000000000001111111111100000000000000000000;
sprite[36] =  50'b00000000000000000000111111111000000000000000000000;
sprite[37] =  50'b00000000000000000000000111000000000000000000000000;
sprite[38] =  50'b00000000000000000000000000000000000000000000000000;
sprite[39] =  50'b00000000000000000000000000000000000000000000000000;
sprite[40] =  50'b00000000000000000000000000000000000000000000000000;
sprite[41] =  50'b00000000000000000000000000000000000000000000000000;
sprite[42] =  50'b00000000000000000000000000000000000000000000000000;
sprite[43] =  50'b00000000000000000000000000000000000000000000000000;
sprite[44] =  50'b00000000000000000000000000000000000000000000000000;
sprite[45] =  50'b00000000000000000000000000000000000000000000000000;
sprite[46] =  50'b00000000000000000000000000000000000000000000000000;
sprite[47] =  50'b00000000000000000000000000000000000000000000000000;
sprite[48] =  50'b00000000000000000000000000000000000000000000000000;
sprite[49] =  50'b00000000000000000000000000000000000000000000000000;
		
		end
		
		4'd6: begin
sprite[0] =  50'b00000000000000000000000000000000000000000000000000;
sprite[1] =  50'b00000000000000000000000000000000000000000000000000;
sprite[2] =  50'b00000000000000000000000000000000000000000000000000;
sprite[3] =  50'b00000000000000000000000000000000000000000000000000;
sprite[4] =  50'b00000000000000000000000000000000000000000000000000;
sprite[5] =  50'b00000000000000000000000000000000000000000000000000;
sprite[6] =  50'b00000000000000000000000000000000000000000000000000;
sprite[7] =  50'b00000000000000000000000000000000000000000000000000;
sprite[8] =  50'b00000000000000000000000000000000000000000000000000;
sprite[9] =  50'b00000000000000000000000000000000000000000000000000;
sprite[10] =  50'b00000000000000000000000000000000000000000000000000;
sprite[11] =  50'b00000000000000000000000000000000000000000000000000;
sprite[12] =  50'b00000000000000000000000000000000000000000000000000;
sprite[13] =  50'b00000000000000000000000001110000000000000000000000;
sprite[14] =  50'b00000000000000000000001111111110000000000000000000;
sprite[15] =  50'b00000000000000000000011111111110000000000000000000;
sprite[16] =  50'b00000000000000000000111100000000000000000000000000;
sprite[17] =  50'b00000000000000000001111000000000000000000000000000;
sprite[18] =  50'b00000000000000000001110000000000000000000000000000;
sprite[19] =  50'b00000000000000000001110000000000000000000000000000;
sprite[20] =  50'b00000000000000000011100000000000000000000000000000;
sprite[21] =  50'b00000000000000000011100000000000000000000000000000;
sprite[22] =  50'b00000000000000000011100011100000000000000000000000;
sprite[23] =  50'b00000000000000000011111111111100000000000000000000;
sprite[24] =  50'b00000000000000000011111111111110000000000000000000;
sprite[25] =  50'b00000000000000000011110000001111000000000000000000;
sprite[26] =  50'b00000000000000000011100000000111000000000000000000;
sprite[27] =  50'b00000000000000000011100000000111000000000000000000;
sprite[28] =  50'b00000000000000000011100000000111000000000000000000;
sprite[29] =  50'b00000000000000000011100000000111000000000000000000;
sprite[30] =  50'b00000000000000000011100000000111000000000000000000;
sprite[31] =  50'b00000000000000000011100000000111000000000000000000;
sprite[32] =  50'b00000000000000000001110000001111000000000000000000;
sprite[33] =  50'b00000000000000000001111000011110000000000000000000;
sprite[34] =  50'b00000000000000000000111111111100000000000000000000;
sprite[35] =  50'b00000000000000000000011111111000000000000000000000;
sprite[36] =  50'b00000000000000000000000011000000000000000000000000;
sprite[37] =  50'b00000000000000000000000000000000000000000000000000;
sprite[38] =  50'b00000000000000000000000000000000000000000000000000;
sprite[39] =  50'b00000000000000000000000000000000000000000000000000;
sprite[40] =  50'b00000000000000000000000000000000000000000000000000;
sprite[41] =  50'b00000000000000000000000000000000000000000000000000;
sprite[42] =  50'b00000000000000000000000000000000000000000000000000;
sprite[43] =  50'b00000000000000000000000000000000000000000000000000;
sprite[44] =  50'b00000000000000000000000000000000000000000000000000;
sprite[45] =  50'b00000000000000000000000000000000000000000000000000;
sprite[46] =  50'b00000000000000000000000000000000000000000000000000;
sprite[47] =  50'b00000000000000000000000000000000000000000000000000;
sprite[48] =  50'b00000000000000000000000000000000000000000000000000;
sprite[49] =  50'b00000000000000000000000000000000000000000000000000;
		
		end
		
		4'd7: begin
sprite[0] =  50'b00000000000000000000000000000000000000000000000000;
sprite[1] =  50'b00000000000000000000000000000000000000000000000000;
sprite[2] =  50'b00000000000000000000000000000000000000000000000000;
sprite[3] =  50'b00000000000000000000000000000000000000000000000000;
sprite[4] =  50'b00000000000000000000000000000000000000000000000000;
sprite[5] =  50'b00000000000000000000000000000000000000000000000000;
sprite[6] =  50'b00000000000000000000000000000000000000000000000000;
sprite[7] =  50'b00000000000000000000000000000000000000000000000000;
sprite[8] =  50'b00000000000000000000000000000000000000000000000000;
sprite[9] =  50'b00000000000000000000000000000000000000000000000000;
sprite[10] =  50'b00000000000000000000000000000000000000000000000000;
sprite[11] =  50'b00000000000000000000000000000000000000000000000000;
sprite[12] =  50'b00000000000000000000000000000000000000000000000000;
sprite[13] =  50'b00000000000000000000000000000000000000000000000000;
sprite[14] =  50'b00000000000000000000000000000000000000000000000000;
sprite[15] =  50'b00000000000000000001111111111111100000000000000000;
sprite[16] =  50'b00000000000000000011111111111111100000000000000000;
sprite[17] =  50'b00000000000000000001111111111111100000000000000000;
sprite[18] =  50'b00000000000000000000000000000111000000000000000000;
sprite[19] =  50'b00000000000000000000000000000111000000000000000000;
sprite[20] =  50'b00000000000000000000000000001110000000000000000000;
sprite[21] =  50'b00000000000000000000000000001110000000000000000000;
sprite[22] =  50'b00000000000000000000000000011110000000000000000000;
sprite[23] =  50'b00000000000000000000000000011100000000000000000000;
sprite[24] =  50'b00000000000000000000000000111100000000000000000000;
sprite[25] =  50'b00000000000000000000000000111000000000000000000000;
sprite[26] =  50'b00000000000000000000000000111000000000000000000000;
sprite[27] =  50'b00000000000000000000000001110000000000000000000000;
sprite[28] =  50'b00000000000000000000000001110000000000000000000000;
sprite[29] =  50'b00000000000000000000000011110000000000000000000000;
sprite[30] =  50'b00000000000000000000000011100000000000000000000000;
sprite[31] =  50'b00000000000000000000000111100000000000000000000000;
sprite[32] =  50'b00000000000000000000000111000000000000000000000000;
sprite[33] =  50'b00000000000000000000001111000000000000000000000000;
sprite[34] =  50'b00000000000000000000001110000000000000000000000000;
sprite[35] =  50'b00000000000000000000001110000000000000000000000000;
sprite[36] =  50'b00000000000000000000011100000000000000000000000000;
sprite[37] =  50'b00000000000000000000000000000000000000000000000000;
sprite[38] =  50'b00000000000000000000000000000000000000000000000000;
sprite[39] =  50'b00000000000000000000000000000000000000000000000000;
sprite[40] =  50'b00000000000000000000000000000000000000000000000000;
sprite[41] =  50'b00000000000000000000000000000000000000000000000000;
sprite[42] =  50'b00000000000000000000000000000000000000000000000000;
sprite[43] =  50'b00000000000000000000000000000000000000000000000000;
sprite[44] =  50'b00000000000000000000000000000000000000000000000000;
sprite[45] =  50'b00000000000000000000000000000000000000000000000000;
sprite[46] =  50'b00000000000000000000000000000000000000000000000000;
sprite[47] =  50'b00000000000000000000000000000000000000000000000000;
sprite[48] =  50'b00000000000000000000000000000000000000000000000000;
sprite[49] =  50'b00000000000000000000000000000000000000000000000000;
		
		end
		
		4'd8: begin
sprite[0] =  50'b00000000000000000000000000000000000000000000000000;
sprite[1] =  50'b00000000000000000000000000000000000000000000000000;
sprite[2] =  50'b00000000000000000000000000000000000000000000000000;
sprite[3] =  50'b00000000000000000000000000000000000000000000000000;
sprite[4] =  50'b00000000000000000000000000000000000000000000000000;
sprite[5] =  50'b00000000000000000000000000000000000000000000000000;
sprite[6] =  50'b00000000000000000000000000000000000000000000000000;
sprite[7] =  50'b00000000000000000000000000000000000000000000000000;
sprite[8] =  50'b00000000000000000000000000000000000000000000000000;
sprite[9] =  50'b00000000000000000000000000000000000000000000000000;
sprite[10] =  50'b00000000000000000000000000000000000000000000000000;
sprite[11] =  50'b00000000000000000000000000000000000000000000000000;
sprite[12] =  50'b00000000000000000000000000000000000000000000000000;
sprite[13] =  50'b00000000000000000000000000000000000000000000000000;
sprite[14] =  50'b00000000000000000000000011100000000000000000000000;
sprite[15] =  50'b00000000000000000000011111111100000000000000000000;
sprite[16] =  50'b00000000000000000000111111111110000000000000000000;
sprite[17] =  50'b00000000000000000000111000001111000000000000000000;
sprite[18] =  50'b00000000000000000001110000000111000000000000000000;
sprite[19] =  50'b00000000000000000001110000000111000000000000000000;
sprite[20] =  50'b00000000000000000001110000000111000000000000000000;
sprite[21] =  50'b00000000000000000001110000000111000000000000000000;
sprite[22] =  50'b00000000000000000000111000001110000000000000000000;
sprite[23] =  50'b00000000000000000000111100011110000000000000000000;
sprite[24] =  50'b00000000000000000000011111111100000000000000000000;
sprite[25] =  50'b00000000000000000000000111111000000000000000000000;
sprite[26] =  50'b00000000000000000000001111111100000000000000000000;
sprite[27] =  50'b00000000000000000000111100111110000000000000000000;
sprite[28] =  50'b00000000000000000001111000001111000000000000000000;
sprite[29] =  50'b00000000000000000001110000000111100000000000000000;
sprite[30] =  50'b00000000000000000011110000000011100000000000000000;
sprite[31] =  50'b00000000000000000011100000000011100000000000000000;
sprite[32] =  50'b00000000000000000011100000000011100000000000000000;
sprite[33] =  50'b00000000000000000011110000000111100000000000000000;
sprite[34] =  50'b00000000000000000001111000001111000000000000000000;
sprite[35] =  50'b00000000000000000000111111111110000000000000000000;
sprite[36] =  50'b00000000000000000000011111111100000000000000000000;
sprite[37] =  50'b00000000000000000000000011100000000000000000000000;
sprite[38] =  50'b00000000000000000000000000000000000000000000000000;
sprite[39] =  50'b00000000000000000000000000000000000000000000000000;
sprite[40] =  50'b00000000000000000000000000000000000000000000000000;
sprite[41] =  50'b00000000000000000000000000000000000000000000000000;
sprite[42] =  50'b00000000000000000000000000000000000000000000000000;
sprite[43] =  50'b00000000000000000000000000000000000000000000000000;
sprite[44] =  50'b00000000000000000000000000000000000000000000000000;
sprite[45] =  50'b00000000000000000000000000000000000000000000000000;
sprite[46] =  50'b00000000000000000000000000000000000000000000000000;
sprite[47] =  50'b00000000000000000000000000000000000000000000000000;
sprite[48] =  50'b00000000000000000000000000000000000000000000000000;
sprite[49] =  50'b00000000000000000000000000000000000000000000000000;
		
		end
		
		4'd9: begin
sprite[0] =  50'b00000000000000000000000000000000000000000000000000;
sprite[1] =  50'b00000000000000000000000000000000000000000000000000;
sprite[2] =  50'b00000000000000000000000000000000000000000000000000;
sprite[3] =  50'b00000000000000000000000000000000000000000000000000;
sprite[4] =  50'b00000000000000000000000000000000000000000000000000;
sprite[5] =  50'b00000000000000000000000000000000000000000000000000;
sprite[6] =  50'b00000000000000000000000000000000000000000000000000;
sprite[7] =  50'b00000000000000000000000000000000000000000000000000;
sprite[8] =  50'b00000000000000000000000000000000000000000000000000;
sprite[9] =  50'b00000000000000000000000000000000000000000000000000;
sprite[10] =  50'b00000000000000000000000000000000000000000000000000;
sprite[11] =  50'b00000000000000000000000000000000000000000000000000;
sprite[12] =  50'b00000000000000000000000011100000000000000000000000;
sprite[13] =  50'b00000000000000000000011111111000000000000000000000;
sprite[14] =  50'b00000000000000000000111111111100000000000000000000;
sprite[15] =  50'b00000000000000000001111000001110000000000000000000;
sprite[16] =  50'b00000000000000000001110000001111000000000000000000;
sprite[17] =  50'b00000000000000000011110000000111000000000000000000;
sprite[18] =  50'b00000000000000000011100000000111000000000000000000;
sprite[19] =  50'b00000000000000000011100000000111000000000000000000;
sprite[20] =  50'b00000000000000000011100000000111100000000000000000;
sprite[21] =  50'b00000000000000000011100000000011100000000000000000;
sprite[22] =  50'b00000000000000000001110000000011100000000000000000;
sprite[23] =  50'b00000000000000000001111000001111100000000000000000;
sprite[24] =  50'b00000000000000000000111111111111100000000000000000;
sprite[25] =  50'b00000000000000000000011111111111100000000000000000;
sprite[26] =  50'b00000000000000000000000011000011000000000000000000;
sprite[27] =  50'b00000000000000000000000000000111000000000000000000;
sprite[28] =  50'b00000000000000000000000000000111000000000000000000;
sprite[29] =  50'b00000000000000000000000000000111000000000000000000;
sprite[30] =  50'b00000000000000000000000000001110000000000000000000;
sprite[31] =  50'b00000000000000000000000000001110000000000000000000;
sprite[32] =  50'b00000000000000000001000000111100000000000000000000;
sprite[33] =  50'b00000000000000000001111111111000000000000000000000;
sprite[34] =  50'b00000000000000000001111111110000000000000000000000;
sprite[35] =  50'b00000000000000000000001110000000000000000000000000;
sprite[36] =  50'b00000000000000000000000000000000000000000000000000;
sprite[37] =  50'b00000000000000000000000000000000000000000000000000;
sprite[38] =  50'b00000000000000000000000000000000000000000000000000;
sprite[39] =  50'b00000000000000000000000000000000000000000000000000;
sprite[40] =  50'b00000000000000000000000000000000000000000000000000;
sprite[41] =  50'b00000000000000000000000000000000000000000000000000;
sprite[42] =  50'b00000000000000000000000000000000000000000000000000;
sprite[43] =  50'b00000000000000000000000000000000000000000000000000;
sprite[44] =  50'b00000000000000000000000000000000000000000000000000;
sprite[45] =  50'b00000000000000000000000000000000000000000000000000;
sprite[46] =  50'b00000000000000000000000000000000000000000000000000;
sprite[47] =  50'b00000000000000000000000000000000000000000000000000;
sprite[48] =  50'b00000000000000000000000000000000000000000000000000;
sprite[49] =  50'b00000000000000000000000000000000000000000000000000;
		
		end
	
	endcase

end 

    wire signed [9:0] x_rel, y_rel;
    assign x_rel = hsync - 505;
    assign y_rel = vsync - 189;
	 
    always @(*) begin
        // Default color is black
        rgb = 24'h000000;
        // Check if the current pixel is within the bounds of the sprite
        if (x_rel >= -25 && x_rel < 25 && y_rel >= -25 && y_rel < 25) begin
            if (sprite[y_rel + 25][x_rel + 25]) begin
                rgb = 24'hFFFF00; 
            end
				else begin
					 rgb=24'h000000;
				end
        end
    end
endmodule